module SumModule(input [31:0] num1, num2, output signed [31:0] result);
    assign result = num1 + num2;
endmodule
